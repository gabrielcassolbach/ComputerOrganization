-- Control Unit