library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity processor is
   port();
end entity;

architecture struct of processor is 

end architecture;